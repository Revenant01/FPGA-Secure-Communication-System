
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ENC_addKey IS

    GENERIC (index : INTEGER);

    PORT (
        inval : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
        outval : OUT STD_LOGIC_VECTOR (127 DOWNTO 0));
END ENC_addKey;

ARCHITECTURE Behavioral OF ENC_addKey IS

    --a088232afa54a36cfe2c397617b13905
    CONSTANT key : STD_LOGIC_VECTOR(1407 DOWNTO 0) := X"2b28ab097eaef7cf15d2154f16a6883ca088232afa54a36cfe2c397617b13905f27a5973c296355995b980f6f2437a7f3d471e6d8016237a47fe7e887d3e443befa8b6db4452710ba55b25ad417f3b00d47cca11d183f2f9c69db815f887bcbc6d11dbca880bf900a33e86937afd41fd4e5f844e545fa6a6f7c94fdc0ef3b24feab5317fd28d2b8d73baf52921d2602fac192867775ad15c66dc2900f321416ed0c9e1b614ee3f63f9250c0ca889c8a6";

BEGIN

    outval <= inval XOR key(index DOWNTO index - 127);

END Behavioral;