LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ENC_SBOX IS
    PORT (
        inval : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        outval : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENC_SBOX;

ARCHITECTURE Behavioral OF ENC_SBOX IS
BEGIN

    PROCESS (inval)
    BEGIN
        CASE inval IS
            WHEN x"00" => outval <= x"63";
            WHEN x"01" => outval <= x"7c";
            WHEN x"02" => outval <= x"77";
            WHEN x"03" => outval <= x"7b";
            WHEN x"04" => outval <= x"f2";
            WHEN x"05" => outval <= x"6b";
            WHEN x"06" => outval <= x"6f";
            WHEN x"07" => outval <= x"c5";
            WHEN x"08" => outval <= x"30";
            WHEN x"09" => outval <= x"01";
            WHEN x"0a" => outval <= x"67";
            WHEN x"0b" => outval <= x"2b";
            WHEN x"0c" => outval <= x"fe";
            WHEN x"0d" => outval <= x"d7";
            WHEN x"0e" => outval <= x"ab";
            WHEN x"0f" => outval <= x"76";
            WHEN x"10" => outval <= x"ca";
            WHEN x"11" => outval <= x"82";
            WHEN x"12" => outval <= x"c9";
            WHEN x"13" => outval <= x"7d";
            WHEN x"14" => outval <= x"fa";
            WHEN x"15" => outval <= x"59";
            WHEN x"16" => outval <= x"47";
            WHEN x"17" => outval <= x"f0";
            WHEN x"18" => outval <= x"ad";
            WHEN x"19" => outval <= x"d4";
            WHEN x"1a" => outval <= x"a2";
            WHEN x"1b" => outval <= x"af";
            WHEN x"1c" => outval <= x"9c";
            WHEN x"1d" => outval <= x"a4";
            WHEN x"1e" => outval <= x"72";
            WHEN x"1f" => outval <= x"c0";
            WHEN x"20" => outval <= x"b7";
            WHEN x"21" => outval <= x"fd";
            WHEN x"22" => outval <= x"93";
            WHEN x"23" => outval <= x"26";
            WHEN x"24" => outval <= x"36";
            WHEN x"25" => outval <= x"3f";
            WHEN x"26" => outval <= x"f7";
            WHEN x"27" => outval <= x"cc";
            WHEN x"28" => outval <= x"34";
            WHEN x"29" => outval <= x"a5";
            WHEN x"2a" => outval <= x"e5";
            WHEN x"2b" => outval <= x"f1";
            WHEN x"2c" => outval <= x"71";
            WHEN x"2d" => outval <= x"d8";
            WHEN x"2e" => outval <= x"31";
            WHEN x"2f" => outval <= x"15";
            WHEN x"30" => outval <= x"04";
            WHEN x"31" => outval <= x"c7";
            WHEN x"32" => outval <= x"23";
            WHEN x"33" => outval <= x"c3";
            WHEN x"34" => outval <= x"18";
            WHEN x"35" => outval <= x"96";
            WHEN x"36" => outval <= x"05";
            WHEN x"37" => outval <= x"9a";
            WHEN x"38" => outval <= x"07";
            WHEN x"39" => outval <= x"12";
            WHEN x"3a" => outval <= x"80";
            WHEN x"3b" => outval <= x"e2";
            WHEN x"3c" => outval <= x"eb";
            WHEN x"3d" => outval <= x"27";
            WHEN x"3e" => outval <= x"b2";
            WHEN x"3f" => outval <= x"75";
            WHEN x"40" => outval <= x"09";
            WHEN x"41" => outval <= x"83";
            WHEN x"42" => outval <= x"2c";
            WHEN x"43" => outval <= x"1a";
            WHEN x"44" => outval <= x"1b";
            WHEN x"45" => outval <= x"6e";
            WHEN x"46" => outval <= x"5a";
            WHEN x"47" => outval <= x"a0";
            WHEN x"48" => outval <= x"52";
            WHEN x"49" => outval <= x"3b";
            WHEN x"4a" => outval <= x"d6";
            WHEN x"4b" => outval <= x"b3";
            WHEN x"4c" => outval <= x"29";
            WHEN x"4d" => outval <= x"e3";
            WHEN x"4e" => outval <= x"2f";
            WHEN x"4f" => outval <= x"84";
            WHEN x"50" => outval <= x"53";
            WHEN x"51" => outval <= x"d1";
            WHEN x"52" => outval <= x"00";
            WHEN x"53" => outval <= x"ed";
            WHEN x"54" => outval <= x"20";
            WHEN x"55" => outval <= x"fc";
            WHEN x"56" => outval <= x"b1";
            WHEN x"57" => outval <= x"5b";
            WHEN x"58" => outval <= x"6a";
            WHEN x"59" => outval <= x"cb";
            WHEN x"5a" => outval <= x"be";
            WHEN x"5b" => outval <= x"39";
            WHEN x"5c" => outval <= x"4a";
            WHEN x"5d" => outval <= x"4c";
            WHEN x"5e" => outval <= x"58";
            WHEN x"5f" => outval <= x"cf";
            WHEN x"60" => outval <= x"d0";
            WHEN x"61" => outval <= x"ef";
            WHEN x"62" => outval <= x"aa";
            WHEN x"63" => outval <= x"fb";
            WHEN x"64" => outval <= x"43";
            WHEN x"65" => outval <= x"4d";
            WHEN x"66" => outval <= x"33";
            WHEN x"67" => outval <= x"85";
            WHEN x"68" => outval <= x"45";
            WHEN x"69" => outval <= x"f9";
            WHEN x"6a" => outval <= x"02";
            WHEN x"6b" => outval <= x"7f";
            WHEN x"6c" => outval <= x"50";
            WHEN x"6d" => outval <= x"3c";
            WHEN x"6e" => outval <= x"9f";
            WHEN x"6f" => outval <= x"a8";
            WHEN x"70" => outval <= x"51";
            WHEN x"71" => outval <= x"a3";
            WHEN x"72" => outval <= x"40";
            WHEN x"73" => outval <= x"8f";
            WHEN x"74" => outval <= x"92";
            WHEN x"75" => outval <= x"9d";
            WHEN x"76" => outval <= x"38";
            WHEN x"77" => outval <= x"f5";
            WHEN x"78" => outval <= x"bc";
            WHEN x"79" => outval <= x"b6";
            WHEN x"7a" => outval <= x"da";
            WHEN x"7b" => outval <= x"21";
            WHEN x"7c" => outval <= x"10";
            WHEN x"7d" => outval <= x"ff";
            WHEN x"7e" => outval <= x"f3";
            WHEN x"7f" => outval <= x"d2";
            WHEN x"80" => outval <= x"cd";
            WHEN x"81" => outval <= x"0c";
            WHEN x"82" => outval <= x"13";
            WHEN x"83" => outval <= x"ec";
            WHEN x"84" => outval <= x"5f";
            WHEN x"85" => outval <= x"97";
            WHEN x"86" => outval <= x"44";
            WHEN x"87" => outval <= x"17";
            WHEN x"88" => outval <= x"c4";
            WHEN x"89" => outval <= x"a7";
            WHEN x"8a" => outval <= x"7e";
            WHEN x"8b" => outval <= x"3d";
            WHEN x"8c" => outval <= x"64";
            WHEN x"8d" => outval <= x"5d";
            WHEN x"8e" => outval <= x"19";
            WHEN x"8f" => outval <= x"73";
            WHEN x"90" => outval <= x"60";
            WHEN x"91" => outval <= x"81";
            WHEN x"92" => outval <= x"4f";
            WHEN x"93" => outval <= x"dc";
            WHEN x"94" => outval <= x"22";
            WHEN x"95" => outval <= x"2a";
            WHEN x"96" => outval <= x"90";
            WHEN x"97" => outval <= x"88";
            WHEN x"98" => outval <= x"46";
            WHEN x"99" => outval <= x"ee";
            WHEN x"9a" => outval <= x"b8";
            WHEN x"9b" => outval <= x"14";
            WHEN x"9c" => outval <= x"de";
            WHEN x"9d" => outval <= x"5e";
            WHEN x"9e" => outval <= x"0b";
            WHEN x"9f" => outval <= x"db";
            WHEN x"a0" => outval <= x"e0";
            WHEN x"a1" => outval <= x"32";
            WHEN x"a2" => outval <= x"3a";
            WHEN x"a3" => outval <= x"0a";
            WHEN x"a4" => outval <= x"49";
            WHEN x"a5" => outval <= x"06";
            WHEN x"a6" => outval <= x"24";
            WHEN x"a7" => outval <= x"5c";
            WHEN x"a8" => outval <= x"c2";
            WHEN x"a9" => outval <= x"d3";
            WHEN x"aa" => outval <= x"ac";
            WHEN x"ab" => outval <= x"62";
            WHEN x"ac" => outval <= x"91";
            WHEN x"ad" => outval <= x"95";
            WHEN x"ae" => outval <= x"e4";
            WHEN x"af" => outval <= x"79";
            WHEN x"b0" => outval <= x"e7";
            WHEN x"b1" => outval <= x"c8";
            WHEN x"b2" => outval <= x"37";
            WHEN x"b3" => outval <= x"6d";
            WHEN x"b4" => outval <= x"8d";
            WHEN x"b5" => outval <= x"d5";
            WHEN x"b6" => outval <= x"4e";
            WHEN x"b7" => outval <= x"a9";
            WHEN x"b8" => outval <= x"6c";
            WHEN x"b9" => outval <= x"56";
            WHEN x"ba" => outval <= x"f4";
            WHEN x"bb" => outval <= x"ea";
            WHEN x"bc" => outval <= x"65";
            WHEN x"bd" => outval <= x"7a";
            WHEN x"be" => outval <= x"ae";
            WHEN x"bf" => outval <= x"08";
            WHEN x"c0" => outval <= x"ba";
            WHEN x"c1" => outval <= x"78";
            WHEN x"c2" => outval <= x"25";
            WHEN x"c3" => outval <= x"2e";
            WHEN x"c4" => outval <= x"1c";
            WHEN x"c5" => outval <= x"a6";
            WHEN x"c6" => outval <= x"b4";
            WHEN x"c7" => outval <= x"c6";
            WHEN x"c8" => outval <= x"e8";
            WHEN x"c9" => outval <= x"dd";
            WHEN x"ca" => outval <= x"74";
            WHEN x"cb" => outval <= x"1f";
            WHEN x"cc" => outval <= x"4b";
            WHEN x"cd" => outval <= x"bd";
            WHEN x"ce" => outval <= x"8b";
            WHEN x"cf" => outval <= x"8a";
            WHEN x"d0" => outval <= x"70";
            WHEN x"d1" => outval <= x"3e";
            WHEN x"d2" => outval <= x"b5";
            WHEN x"d3" => outval <= x"66";
            WHEN x"d4" => outval <= x"48";
            WHEN x"d5" => outval <= x"03";
            WHEN x"d6" => outval <= x"f6";
            WHEN x"d7" => outval <= x"0e";
            WHEN x"d8" => outval <= x"61";
            WHEN x"d9" => outval <= x"35";
            WHEN x"da" => outval <= x"57";
            WHEN x"db" => outval <= x"b9";
            WHEN x"dc" => outval <= x"86";
            WHEN x"dd" => outval <= x"c1";
            WHEN x"de" => outval <= x"1d";
            WHEN x"df" => outval <= x"9e";
            WHEN x"e0" => outval <= x"e1";
            WHEN x"e1" => outval <= x"f8";
            WHEN x"e2" => outval <= x"98";
            WHEN x"e3" => outval <= x"11";
            WHEN x"e4" => outval <= x"69";
            WHEN x"e5" => outval <= x"d9";
            WHEN x"e6" => outval <= x"8e";
            WHEN x"e7" => outval <= x"94";
            WHEN x"e8" => outval <= x"9b";
            WHEN x"e9" => outval <= x"1e";
            WHEN x"ea" => outval <= x"87";
            WHEN x"eb" => outval <= x"e9";
            WHEN x"ec" => outval <= x"ce";
            WHEN x"ed" => outval <= x"55";
            WHEN x"ee" => outval <= x"28";
            WHEN x"ef" => outval <= x"df";
            WHEN x"f0" => outval <= x"8c";
            WHEN x"f1" => outval <= x"a1";
            WHEN x"f2" => outval <= x"89";
            WHEN x"f3" => outval <= x"0d";
            WHEN x"f4" => outval <= x"bf";
            WHEN x"f5" => outval <= x"e6";
            WHEN x"f6" => outval <= x"42";
            WHEN x"f7" => outval <= x"68";
            WHEN x"f8" => outval <= x"41";
            WHEN x"f9" => outval <= x"99";
            WHEN x"fa" => outval <= x"2d";
            WHEN x"fb" => outval <= x"0f";
            WHEN x"fc" => outval <= x"b0";
            WHEN x"fd" => outval <= x"54";
            WHEN x"fe" => outval <= x"bb";
            WHEN x"ff" => outval <= x"16";
            WHEN OTHERS => NULL; -- GHDL complains without this statement
        END CASE;

    END PROCESS;
END Behavioral;